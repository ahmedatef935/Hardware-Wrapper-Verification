echo
echo "!!! Pre run"

help

run

echo "!!! Post run"

exec urg -help
exec urg -dir simv.vdb

echo "!!! Post urg"
echo
